 
 


typedef struct packed {
    logic cosim_stop;
    logic cosim_val;
    logic cosim_go; 
    logic cosim_done; 
    
 } control;